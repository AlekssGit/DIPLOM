library verilog;
use verilog.vl_types.all;
entity SPI_vlg_vec_tst is
end SPI_vlg_vec_tst;
